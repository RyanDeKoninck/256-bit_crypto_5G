//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Ryan De Koninck
// 
// Create Date: 04/20/2023 15:12:00
// Design Name: 
// Module Name: zuc256_sbox1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`default_nettype none

module zuc256_sbox(
                input wire [31 : 0]  sboxw,
                output wire [31 : 0] new_sboxw
               );


  //----------------------------------------------------------------
  // The sbox array.
  //----------------------------------------------------------------
  wire [7 : 0] sbox0 [0 : 255];
  wire [7 : 0] sbox1 [0 : 255];


  //----------------------------------------------------------------
  // Four parallel muxes.
  //----------------------------------------------------------------
  assign new_sboxw[31 : 24] = sbox0[sboxw[31 : 24]];
  assign new_sboxw[23 : 16] = sbox1[sboxw[23 : 16]];
  assign new_sboxw[15 : 08] = sbox0[sboxw[15 : 08]];
  assign new_sboxw[07 : 00] = sbox1[sboxw[07 : 00]];


  //----------------------------------------------------------------
  // Creating the sbox array contents.
  //----------------------------------------------------------------
   assign sbox0[8'h0] = 8'h3e;
   assign sbox0[8'h1] = 8'h72;
   assign sbox0[8'h2] = 8'h5b;
   assign sbox0[8'h3] = 8'h47;
   assign sbox0[8'h4] = 8'hca;
   assign sbox0[8'h5] = 8'he0;
   assign sbox0[8'h6] = 8'h0;
   assign sbox0[8'h7] = 8'h33;
   assign sbox0[8'h8] = 8'h4;
   assign sbox0[8'h9] = 8'hd1;
   assign sbox0[8'ha] = 8'h54;
   assign sbox0[8'hb] = 8'h98;
   assign sbox0[8'hc] = 8'h9;
   assign sbox0[8'hd] = 8'hb9;
   assign sbox0[8'he] = 8'h6d;
   assign sbox0[8'hf] = 8'hcb;
   assign sbox0[8'h10] = 8'h7b;
   assign sbox0[8'h11] = 8'h1b;
   assign sbox0[8'h12] = 8'hf9;
   assign sbox0[8'h13] = 8'h32;
   assign sbox0[8'h14] = 8'haf;
   assign sbox0[8'h15] = 8'h9d;
   assign sbox0[8'h16] = 8'h6a;
   assign sbox0[8'h17] = 8'ha5;
   assign sbox0[8'h18] = 8'hb8;
   assign sbox0[8'h19] = 8'h2d;
   assign sbox0[8'h1a] = 8'hfc;
   assign sbox0[8'h1b] = 8'h1d;
   assign sbox0[8'h1c] = 8'h8;
   assign sbox0[8'h1d] = 8'h53;
   assign sbox0[8'h1e] = 8'h3;
   assign sbox0[8'h1f] = 8'h90;
   assign sbox0[8'h20] = 8'h4d;
   assign sbox0[8'h21] = 8'h4e;
   assign sbox0[8'h22] = 8'h84;
   assign sbox0[8'h23] = 8'h99;
   assign sbox0[8'h24] = 8'he4;
   assign sbox0[8'h25] = 8'hce;
   assign sbox0[8'h26] = 8'hd9;
   assign sbox0[8'h27] = 8'h91;
   assign sbox0[8'h28] = 8'hdd;
   assign sbox0[8'h29] = 8'hb6;
   assign sbox0[8'h2a] = 8'h85;
   assign sbox0[8'h2b] = 8'h48;
   assign sbox0[8'h2c] = 8'h8b;
   assign sbox0[8'h2d] = 8'h29;
   assign sbox0[8'h2e] = 8'h6e;
   assign sbox0[8'h2f] = 8'hac;
   assign sbox0[8'h30] = 8'hcd;
   assign sbox0[8'h31] = 8'hc1;
   assign sbox0[8'h32] = 8'hf8;
   assign sbox0[8'h33] = 8'h1e;
   assign sbox0[8'h34] = 8'h73;
   assign sbox0[8'h35] = 8'h43;
   assign sbox0[8'h36] = 8'h69;
   assign sbox0[8'h37] = 8'hc6;
   assign sbox0[8'h38] = 8'hb5;
   assign sbox0[8'h39] = 8'hbd;
   assign sbox0[8'h3a] = 8'hfd;
   assign sbox0[8'h3b] = 8'h39;
   assign sbox0[8'h3c] = 8'h63;
   assign sbox0[8'h3d] = 8'h20;
   assign sbox0[8'h3e] = 8'hd4;
   assign sbox0[8'h3f] = 8'h38;
   assign sbox0[8'h40] = 8'h76;
   assign sbox0[8'h41] = 8'h7d;
   assign sbox0[8'h42] = 8'hb2;
   assign sbox0[8'h43] = 8'ha7;
   assign sbox0[8'h44] = 8'hcf;
   assign sbox0[8'h45] = 8'hed;
   assign sbox0[8'h46] = 8'h57;
   assign sbox0[8'h47] = 8'hc5;
   assign sbox0[8'h48] = 8'hf3;
   assign sbox0[8'h49] = 8'h2c;
   assign sbox0[8'h4a] = 8'hbb;
   assign sbox0[8'h4b] = 8'h14;
   assign sbox0[8'h4c] = 8'h21;
   assign sbox0[8'h4d] = 8'h6;
   assign sbox0[8'h4e] = 8'h55;
   assign sbox0[8'h4f] = 8'h9b;
   assign sbox0[8'h50] = 8'he3;
   assign sbox0[8'h51] = 8'hef;
   assign sbox0[8'h52] = 8'h5e;
   assign sbox0[8'h53] = 8'h31;
   assign sbox0[8'h54] = 8'h4f;
   assign sbox0[8'h55] = 8'h7f;
   assign sbox0[8'h56] = 8'h5a;
   assign sbox0[8'h57] = 8'ha4;
   assign sbox0[8'h58] = 8'hd;
   assign sbox0[8'h59] = 8'h82;
   assign sbox0[8'h5a] = 8'h51;
   assign sbox0[8'h5b] = 8'h49;
   assign sbox0[8'h5c] = 8'h5f;
   assign sbox0[8'h5d] = 8'hba;
   assign sbox0[8'h5e] = 8'h58;
   assign sbox0[8'h5f] = 8'h1c;
   assign sbox0[8'h60] = 8'h4a;
   assign sbox0[8'h61] = 8'h16;
   assign sbox0[8'h62] = 8'hd5;
   assign sbox0[8'h63] = 8'h17;
   assign sbox0[8'h64] = 8'ha8;
   assign sbox0[8'h65] = 8'h92;
   assign sbox0[8'h66] = 8'h24;
   assign sbox0[8'h67] = 8'h1f;
   assign sbox0[8'h68] = 8'h8c;
   assign sbox0[8'h69] = 8'hff;
   assign sbox0[8'h6a] = 8'hd8;
   assign sbox0[8'h6b] = 8'hae;
   assign sbox0[8'h6c] = 8'h2e;
   assign sbox0[8'h6d] = 8'h1;
   assign sbox0[8'h6e] = 8'hd3;
   assign sbox0[8'h6f] = 8'had;
   assign sbox0[8'h70] = 8'h3b;
   assign sbox0[8'h71] = 8'h4b;
   assign sbox0[8'h72] = 8'hda;
   assign sbox0[8'h73] = 8'h46;
   assign sbox0[8'h74] = 8'heb;
   assign sbox0[8'h75] = 8'hc9;
   assign sbox0[8'h76] = 8'hde;
   assign sbox0[8'h77] = 8'h9a;
   assign sbox0[8'h78] = 8'h8f;
   assign sbox0[8'h79] = 8'h87;
   assign sbox0[8'h7a] = 8'hd7;
   assign sbox0[8'h7b] = 8'h3a;
   assign sbox0[8'h7c] = 8'h80;
   assign sbox0[8'h7d] = 8'h6f;
   assign sbox0[8'h7e] = 8'h2f;
   assign sbox0[8'h7f] = 8'hc8;
   assign sbox0[8'h80] = 8'hb1;
   assign sbox0[8'h81] = 8'hb4;
   assign sbox0[8'h82] = 8'h37;
   assign sbox0[8'h83] = 8'hf7;
   assign sbox0[8'h84] = 8'ha;
   assign sbox0[8'h85] = 8'h22;
   assign sbox0[8'h86] = 8'h13;
   assign sbox0[8'h87] = 8'h28;
   assign sbox0[8'h88] = 8'h7c;
   assign sbox0[8'h89] = 8'hcc;
   assign sbox0[8'h8a] = 8'h3c;
   assign sbox0[8'h8b] = 8'h89;
   assign sbox0[8'h8c] = 8'hc7;
   assign sbox0[8'h8d] = 8'hc3;
   assign sbox0[8'h8e] = 8'h96;
   assign sbox0[8'h8f] = 8'h56;
   assign sbox0[8'h90] = 8'h7;
   assign sbox0[8'h91] = 8'hbf;
   assign sbox0[8'h92] = 8'h7e;
   assign sbox0[8'h93] = 8'hf0;
   assign sbox0[8'h94] = 8'hb;
   assign sbox0[8'h95] = 8'h2b;
   assign sbox0[8'h96] = 8'h97;
   assign sbox0[8'h97] = 8'h52;
   assign sbox0[8'h98] = 8'h35;
   assign sbox0[8'h99] = 8'h41;
   assign sbox0[8'h9a] = 8'h79;
   assign sbox0[8'h9b] = 8'h61;
   assign sbox0[8'h9c] = 8'ha6;
   assign sbox0[8'h9d] = 8'h4c;
   assign sbox0[8'h9e] = 8'h10;
   assign sbox0[8'h9f] = 8'hfe;
   assign sbox0[8'ha0] = 8'hbc;
   assign sbox0[8'ha1] = 8'h26;
   assign sbox0[8'ha2] = 8'h95;
   assign sbox0[8'ha3] = 8'h88;
   assign sbox0[8'ha4] = 8'h8a;
   assign sbox0[8'ha5] = 8'hb0;
   assign sbox0[8'ha6] = 8'ha3;
   assign sbox0[8'ha7] = 8'hfb;
   assign sbox0[8'ha8] = 8'hc0;
   assign sbox0[8'ha9] = 8'h18;
   assign sbox0[8'haa] = 8'h94;
   assign sbox0[8'hab] = 8'hf2;
   assign sbox0[8'hac] = 8'he1;
   assign sbox0[8'had] = 8'he5;
   assign sbox0[8'hae] = 8'he9;
   assign sbox0[8'haf] = 8'h5d;
   assign sbox0[8'hb0] = 8'hd0;
   assign sbox0[8'hb1] = 8'hdc;
   assign sbox0[8'hb2] = 8'h11;
   assign sbox0[8'hb3] = 8'h66;
   assign sbox0[8'hb4] = 8'h64;
   assign sbox0[8'hb5] = 8'h5c;
   assign sbox0[8'hb6] = 8'hec;
   assign sbox0[8'hb7] = 8'h59;
   assign sbox0[8'hb8] = 8'h42;
   assign sbox0[8'hb9] = 8'h75;
   assign sbox0[8'hba] = 8'h12;
   assign sbox0[8'hbb] = 8'hf5;
   assign sbox0[8'hbc] = 8'h74;
   assign sbox0[8'hbd] = 8'h9c;
   assign sbox0[8'hbe] = 8'haa;
   assign sbox0[8'hbf] = 8'h23;
   assign sbox0[8'hc0] = 8'he;
   assign sbox0[8'hc1] = 8'h86;
   assign sbox0[8'hc2] = 8'hab;
   assign sbox0[8'hc3] = 8'hbe;
   assign sbox0[8'hc4] = 8'h2a;
   assign sbox0[8'hc5] = 8'h2;
   assign sbox0[8'hc6] = 8'he7;
   assign sbox0[8'hc7] = 8'h67;
   assign sbox0[8'hc8] = 8'he6;
   assign sbox0[8'hc9] = 8'h44;
   assign sbox0[8'hca] = 8'ha2;
   assign sbox0[8'hcb] = 8'h6c;
   assign sbox0[8'hcc] = 8'hc2;
   assign sbox0[8'hcd] = 8'h93;
   assign sbox0[8'hce] = 8'h9f;
   assign sbox0[8'hcf] = 8'hf1;
   assign sbox0[8'hd0] = 8'hf6;
   assign sbox0[8'hd1] = 8'hfa;
   assign sbox0[8'hd2] = 8'h36;
   assign sbox0[8'hd3] = 8'hd2;
   assign sbox0[8'hd4] = 8'h50;
   assign sbox0[8'hd5] = 8'h68;
   assign sbox0[8'hd6] = 8'h9e;
   assign sbox0[8'hd7] = 8'h62;
   assign sbox0[8'hd8] = 8'h71;
   assign sbox0[8'hd9] = 8'h15;
   assign sbox0[8'hda] = 8'h3d;
   assign sbox0[8'hdb] = 8'hd6;
   assign sbox0[8'hdc] = 8'h40;
   assign sbox0[8'hdd] = 8'hc4;
   assign sbox0[8'hde] = 8'he2;
   assign sbox0[8'hdf] = 8'hf;
   assign sbox0[8'he0] = 8'h8e;
   assign sbox0[8'he1] = 8'h83;
   assign sbox0[8'he2] = 8'h77;
   assign sbox0[8'he3] = 8'h6b;
   assign sbox0[8'he4] = 8'h25;
   assign sbox0[8'he5] = 8'h5;
   assign sbox0[8'he6] = 8'h3f;
   assign sbox0[8'he7] = 8'hc;
   assign sbox0[8'he8] = 8'h30;
   assign sbox0[8'he9] = 8'hea;
   assign sbox0[8'hea] = 8'h70;
   assign sbox0[8'heb] = 8'hb7;
   assign sbox0[8'hec] = 8'ha1;
   assign sbox0[8'hed] = 8'he8;
   assign sbox0[8'hee] = 8'ha9;
   assign sbox0[8'hef] = 8'h65;
   assign sbox0[8'hf0] = 8'h8d;
   assign sbox0[8'hf1] = 8'h27;
   assign sbox0[8'hf2] = 8'h1a;
   assign sbox0[8'hf3] = 8'hdb;
   assign sbox0[8'hf4] = 8'h81;
   assign sbox0[8'hf5] = 8'hb3;
   assign sbox0[8'hf6] = 8'ha0;
   assign sbox0[8'hf7] = 8'hf4;
   assign sbox0[8'hf8] = 8'h45;
   assign sbox0[8'hf9] = 8'h7a;
   assign sbox0[8'hfa] = 8'h19;
   assign sbox0[8'hfb] = 8'hdf;
   assign sbox0[8'hfc] = 8'hee;
   assign sbox0[8'hfd] = 8'h78;
   assign sbox0[8'hfe] = 8'h34;
   assign sbox0[8'hff] = 8'h60;
   
   assign sbox1[8'h0] = 8'h55;
   assign sbox1[8'h1] = 8'hc2;
   assign sbox1[8'h2] = 8'h63;
   assign sbox1[8'h3] = 8'h71;
   assign sbox1[8'h4] = 8'h3b;
   assign sbox1[8'h5] = 8'hc8;
   assign sbox1[8'h6] = 8'h47;
   assign sbox1[8'h7] = 8'h86;
   assign sbox1[8'h8] = 8'h9f;
   assign sbox1[8'h9] = 8'h3c;
   assign sbox1[8'ha] = 8'hda;
   assign sbox1[8'hb] = 8'h5b;
   assign sbox1[8'hc] = 8'h29;
   assign sbox1[8'hd] = 8'haa;
   assign sbox1[8'he] = 8'hfd;
   assign sbox1[8'hf] = 8'h77;
   assign sbox1[8'h10] = 8'h8c;
   assign sbox1[8'h11] = 8'hc5;
   assign sbox1[8'h12] = 8'h94;
   assign sbox1[8'h13] = 8'hc;
   assign sbox1[8'h14] = 8'ha6;
   assign sbox1[8'h15] = 8'h1a;
   assign sbox1[8'h16] = 8'h13;
   assign sbox1[8'h17] = 8'h0;
   assign sbox1[8'h18] = 8'he3;
   assign sbox1[8'h19] = 8'ha8;
   assign sbox1[8'h1a] = 8'h16;
   assign sbox1[8'h1b] = 8'h72;
   assign sbox1[8'h1c] = 8'h40;
   assign sbox1[8'h1d] = 8'hf9;
   assign sbox1[8'h1e] = 8'hf8;
   assign sbox1[8'h1f] = 8'h42;
   assign sbox1[8'h20] = 8'h44;
   assign sbox1[8'h21] = 8'h26;
   assign sbox1[8'h22] = 8'h68;
   assign sbox1[8'h23] = 8'h96;
   assign sbox1[8'h24] = 8'h81;
   assign sbox1[8'h25] = 8'hd9;
   assign sbox1[8'h26] = 8'h45;
   assign sbox1[8'h27] = 8'h3e;
   assign sbox1[8'h28] = 8'h10;
   assign sbox1[8'h29] = 8'h76;
   assign sbox1[8'h2a] = 8'hc6;
   assign sbox1[8'h2b] = 8'ha7;
   assign sbox1[8'h2c] = 8'h8b;
   assign sbox1[8'h2d] = 8'h39;
   assign sbox1[8'h2e] = 8'h43;
   assign sbox1[8'h2f] = 8'he1;
   assign sbox1[8'h30] = 8'h3a;
   assign sbox1[8'h31] = 8'hb5;
   assign sbox1[8'h32] = 8'h56;
   assign sbox1[8'h33] = 8'h2a;
   assign sbox1[8'h34] = 8'hc0;
   assign sbox1[8'h35] = 8'h6d;
   assign sbox1[8'h36] = 8'hb3;
   assign sbox1[8'h37] = 8'h5;
   assign sbox1[8'h38] = 8'h22;
   assign sbox1[8'h39] = 8'h66;
   assign sbox1[8'h3a] = 8'hbf;
   assign sbox1[8'h3b] = 8'hdc;
   assign sbox1[8'h3c] = 8'hb;
   assign sbox1[8'h3d] = 8'hfa;
   assign sbox1[8'h3e] = 8'h62;
   assign sbox1[8'h3f] = 8'h48;
   assign sbox1[8'h40] = 8'hdd;
   assign sbox1[8'h41] = 8'h20;
   assign sbox1[8'h42] = 8'h11;
   assign sbox1[8'h43] = 8'h6;
   assign sbox1[8'h44] = 8'h36;
   assign sbox1[8'h45] = 8'hc9;
   assign sbox1[8'h46] = 8'hc1;
   assign sbox1[8'h47] = 8'hcf;
   assign sbox1[8'h48] = 8'hf6;
   assign sbox1[8'h49] = 8'h27;
   assign sbox1[8'h4a] = 8'h52;
   assign sbox1[8'h4b] = 8'hbb;
   assign sbox1[8'h4c] = 8'h69;
   assign sbox1[8'h4d] = 8'hf5;
   assign sbox1[8'h4e] = 8'hd4;
   assign sbox1[8'h4f] = 8'h87;
   assign sbox1[8'h50] = 8'h7f;
   assign sbox1[8'h51] = 8'h84;
   assign sbox1[8'h52] = 8'h4c;
   assign sbox1[8'h53] = 8'hd2;
   assign sbox1[8'h54] = 8'h9c;
   assign sbox1[8'h55] = 8'h57;
   assign sbox1[8'h56] = 8'ha4;
   assign sbox1[8'h57] = 8'hbc;
   assign sbox1[8'h58] = 8'h4f;
   assign sbox1[8'h59] = 8'h9a;
   assign sbox1[8'h5a] = 8'hdf;
   assign sbox1[8'h5b] = 8'hfe;
   assign sbox1[8'h5c] = 8'hd6;
   assign sbox1[8'h5d] = 8'h8d;
   assign sbox1[8'h5e] = 8'h7a;
   assign sbox1[8'h5f] = 8'heb;
   assign sbox1[8'h60] = 8'h2b;
   assign sbox1[8'h61] = 8'h53;
   assign sbox1[8'h62] = 8'hd8;
   assign sbox1[8'h63] = 8'h5c;
   assign sbox1[8'h64] = 8'ha1;
   assign sbox1[8'h65] = 8'h14;
   assign sbox1[8'h66] = 8'h17;
   assign sbox1[8'h67] = 8'hfb;
   assign sbox1[8'h68] = 8'h23;
   assign sbox1[8'h69] = 8'hd5;
   assign sbox1[8'h6a] = 8'h7d;
   assign sbox1[8'h6b] = 8'h30;
   assign sbox1[8'h6c] = 8'h67;
   assign sbox1[8'h6d] = 8'h73;
   assign sbox1[8'h6e] = 8'h8;
   assign sbox1[8'h6f] = 8'h9;
   assign sbox1[8'h70] = 8'hee;
   assign sbox1[8'h71] = 8'hb7;
   assign sbox1[8'h72] = 8'h70;
   assign sbox1[8'h73] = 8'h3f;
   assign sbox1[8'h74] = 8'h61;
   assign sbox1[8'h75] = 8'hb2;
   assign sbox1[8'h76] = 8'h19;
   assign sbox1[8'h77] = 8'h8e;
   assign sbox1[8'h78] = 8'h4e;
   assign sbox1[8'h79] = 8'he5;
   assign sbox1[8'h7a] = 8'h4b;
   assign sbox1[8'h7b] = 8'h93;
   assign sbox1[8'h7c] = 8'h8f;
   assign sbox1[8'h7d] = 8'h5d;
   assign sbox1[8'h7e] = 8'hdb;
   assign sbox1[8'h7f] = 8'ha9;
   assign sbox1[8'h80] = 8'had;
   assign sbox1[8'h81] = 8'hf1;
   assign sbox1[8'h82] = 8'hae;
   assign sbox1[8'h83] = 8'h2e;
   assign sbox1[8'h84] = 8'hcb;
   assign sbox1[8'h85] = 8'hd;
   assign sbox1[8'h86] = 8'hfc;
   assign sbox1[8'h87] = 8'hf4;
   assign sbox1[8'h88] = 8'h2d;
   assign sbox1[8'h89] = 8'h46;
   assign sbox1[8'h8a] = 8'h6e;
   assign sbox1[8'h8b] = 8'h1d;
   assign sbox1[8'h8c] = 8'h97;
   assign sbox1[8'h8d] = 8'he8;
   assign sbox1[8'h8e] = 8'hd1;
   assign sbox1[8'h8f] = 8'he9;
   assign sbox1[8'h90] = 8'h4d;
   assign sbox1[8'h91] = 8'h37;
   assign sbox1[8'h92] = 8'ha5;
   assign sbox1[8'h93] = 8'h75;
   assign sbox1[8'h94] = 8'h5e;
   assign sbox1[8'h95] = 8'h83;
   assign sbox1[8'h96] = 8'h9e;
   assign sbox1[8'h97] = 8'hab;
   assign sbox1[8'h98] = 8'h82;
   assign sbox1[8'h99] = 8'h9d;
   assign sbox1[8'h9a] = 8'hb9;
   assign sbox1[8'h9b] = 8'h1c;
   assign sbox1[8'h9c] = 8'he0;
   assign sbox1[8'h9d] = 8'hcd;
   assign sbox1[8'h9e] = 8'h49;
   assign sbox1[8'h9f] = 8'h89;
   assign sbox1[8'ha0] = 8'h1;
   assign sbox1[8'ha1] = 8'hb6;
   assign sbox1[8'ha2] = 8'hbd;
   assign sbox1[8'ha3] = 8'h58;
   assign sbox1[8'ha4] = 8'h24;
   assign sbox1[8'ha5] = 8'ha2;
   assign sbox1[8'ha6] = 8'h5f;
   assign sbox1[8'ha7] = 8'h38;
   assign sbox1[8'ha8] = 8'h78;
   assign sbox1[8'ha9] = 8'h99;
   assign sbox1[8'haa] = 8'h15;
   assign sbox1[8'hab] = 8'h90;
   assign sbox1[8'hac] = 8'h50;
   assign sbox1[8'had] = 8'hb8;
   assign sbox1[8'hae] = 8'h95;
   assign sbox1[8'haf] = 8'he4;
   assign sbox1[8'hb0] = 8'hd0;
   assign sbox1[8'hb1] = 8'h91;
   assign sbox1[8'hb2] = 8'hc7;
   assign sbox1[8'hb3] = 8'hce;
   assign sbox1[8'hb4] = 8'hed;
   assign sbox1[8'hb5] = 8'hf;
   assign sbox1[8'hb6] = 8'hb4;
   assign sbox1[8'hb7] = 8'h6f;
   assign sbox1[8'hb8] = 8'ha0;
   assign sbox1[8'hb9] = 8'hcc;
   assign sbox1[8'hba] = 8'hf0;
   assign sbox1[8'hbb] = 8'h2;
   assign sbox1[8'hbc] = 8'h4a;
   assign sbox1[8'hbd] = 8'h79;
   assign sbox1[8'hbe] = 8'hc3;
   assign sbox1[8'hbf] = 8'hde;
   assign sbox1[8'hc0] = 8'ha3;
   assign sbox1[8'hc1] = 8'hef;
   assign sbox1[8'hc2] = 8'hea;
   assign sbox1[8'hc3] = 8'h51;
   assign sbox1[8'hc4] = 8'he6;
   assign sbox1[8'hc5] = 8'h6b;
   assign sbox1[8'hc6] = 8'h18;
   assign sbox1[8'hc7] = 8'hec;
   assign sbox1[8'hc8] = 8'h1b;
   assign sbox1[8'hc9] = 8'h2c;
   assign sbox1[8'hca] = 8'h80;
   assign sbox1[8'hcb] = 8'hf7;
   assign sbox1[8'hcc] = 8'h74;
   assign sbox1[8'hcd] = 8'he7;
   assign sbox1[8'hce] = 8'hff;
   assign sbox1[8'hcf] = 8'h21;
   assign sbox1[8'hd0] = 8'h5a;
   assign sbox1[8'hd1] = 8'h6a;
   assign sbox1[8'hd2] = 8'h54;
   assign sbox1[8'hd3] = 8'h1e;
   assign sbox1[8'hd4] = 8'h41;
   assign sbox1[8'hd5] = 8'h31;
   assign sbox1[8'hd6] = 8'h92;
   assign sbox1[8'hd7] = 8'h35;
   assign sbox1[8'hd8] = 8'hc4;
   assign sbox1[8'hd9] = 8'h33;
   assign sbox1[8'hda] = 8'h7;
   assign sbox1[8'hdb] = 8'ha;
   assign sbox1[8'hdc] = 8'hba;
   assign sbox1[8'hdd] = 8'h7e;
   assign sbox1[8'hde] = 8'he;
   assign sbox1[8'hdf] = 8'h34;
   assign sbox1[8'he0] = 8'h88;
   assign sbox1[8'he1] = 8'hb1;
   assign sbox1[8'he2] = 8'h98;
   assign sbox1[8'he3] = 8'h7c;
   assign sbox1[8'he4] = 8'hf3;
   assign sbox1[8'he5] = 8'h3d;
   assign sbox1[8'he6] = 8'h60;
   assign sbox1[8'he7] = 8'h6c;
   assign sbox1[8'he8] = 8'h7b;
   assign sbox1[8'he9] = 8'hca;
   assign sbox1[8'hea] = 8'hd3;
   assign sbox1[8'heb] = 8'h1f;
   assign sbox1[8'hec] = 8'h32;
   assign sbox1[8'hed] = 8'h65;
   assign sbox1[8'hee] = 8'h4;
   assign sbox1[8'hef] = 8'h28;
   assign sbox1[8'hf0] = 8'h64;
   assign sbox1[8'hf1] = 8'hbe;
   assign sbox1[8'hf2] = 8'h85;
   assign sbox1[8'hf3] = 8'h9b;
   assign sbox1[8'hf4] = 8'h2f;
   assign sbox1[8'hf5] = 8'h59;
   assign sbox1[8'hf6] = 8'h8a;
   assign sbox1[8'hf7] = 8'hd7;
   assign sbox1[8'hf8] = 8'hb0;
   assign sbox1[8'hf9] = 8'h25;
   assign sbox1[8'hfa] = 8'hac;
   assign sbox1[8'hfb] = 8'haf;
   assign sbox1[8'hfc] = 8'h12;
   assign sbox1[8'hfd] = 8'h3;
   assign sbox1[8'hfe] = 8'he2;
   assign sbox1[8'hff] = 8'hf2;

endmodule // zuc256_sbox

//======================================================================
// EOF zuc256_sbox.v
//======================================================================
